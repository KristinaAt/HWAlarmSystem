-- Copyright (C) 1991-2011 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 11.1 Build 259 01/25/2012 Service Pack 2 SJ Web Edition"
-- CREATED		"Sun Jan 20 00:44:32 2019"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY dlock IS 
	PORT
	(
		DATA :  IN  STD_LOGIC;
		CLOCK :  IN  STD_LOGIC;
		RESET :  IN  STD_LOGIC;
		LOCK :  OUT  STD_LOGIC;
		ALARM :  OUT  STD_LOGIC
	);
END dlock;

ARCHITECTURE bdf_type OF dlock IS 

SIGNAL	negDATAandNQ2 :  STD_LOGIC;
SIGNAL	NQ0 :  STD_LOGIC;
SIGNAL	NQ1 :  STD_LOGIC;
SIGNAL	NQ2 :  STD_LOGIC;
SIGNAL	Q0 :  STD_LOGIC;
SIGNAL	Q1 :  STD_LOGIC;
SIGNAL	Q2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_2 <= '1';
SYNTHESIZED_WIRE_5 <= '1';
SYNTHESIZED_WIRE_8 <= '1';



PROCESS(CLOCK,SYNTHESIZED_WIRE_22,SYNTHESIZED_WIRE_2)
BEGIN
IF (SYNTHESIZED_WIRE_22 = '0') THEN
	Q2 <= '0';
ELSIF (SYNTHESIZED_WIRE_2 = '0') THEN
	Q2 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	Q2 <= SYNTHESIZED_WIRE_1;
END IF;
END PROCESS;


PROCESS(CLOCK,SYNTHESIZED_WIRE_22,SYNTHESIZED_WIRE_5)
BEGIN
IF (SYNTHESIZED_WIRE_22 = '0') THEN
	Q1 <= '0';
ELSIF (SYNTHESIZED_WIRE_5 = '0') THEN
	Q1 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	Q1 <= SYNTHESIZED_WIRE_4;
END IF;
END PROCESS;



PROCESS(CLOCK,SYNTHESIZED_WIRE_22,SYNTHESIZED_WIRE_8)
BEGIN
IF (SYNTHESIZED_WIRE_22 = '0') THEN
	Q0 <= '0';
ELSIF (SYNTHESIZED_WIRE_8 = '0') THEN
	Q0 <= '1';
ELSIF (RISING_EDGE(CLOCK)) THEN
	Q0 <= SYNTHESIZED_WIRE_7;
END IF;
END PROCESS;




SYNTHESIZED_WIRE_22 <= NOT(RESET);



SYNTHESIZED_WIRE_19 <= NOT(DATA XOR Q2);


SYNTHESIZED_WIRE_7 <= NOT(SYNTHESIZED_WIRE_9 AND SYNTHESIZED_WIRE_10 AND SYNTHESIZED_WIRE_11);


SYNTHESIZED_WIRE_4 <= NOT(NQ0 AND negDATAandNQ2 AND SYNTHESIZED_WIRE_23);


SYNTHESIZED_WIRE_1 <= NOT(SYNTHESIZED_WIRE_13 AND SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_15);


NQ2 <= NOT(Q2);



SYNTHESIZED_WIRE_13 <= NOT(SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17);


SYNTHESIZED_WIRE_15 <= NOT(Q0 AND SYNTHESIZED_WIRE_18);


SYNTHESIZED_WIRE_23 <= NOT(DATA AND NQ1 AND NQ0);


negDATAandNQ2 <= NOT(NQ2 AND DATA);


SYNTHESIZED_WIRE_9 <= NOT(SYNTHESIZED_WIRE_19 AND Q0);


SYNTHESIZED_WIRE_10 <= NOT(NQ0 AND SYNTHESIZED_WIRE_20);


SYNTHESIZED_WIRE_11 <= Q1 XOR Q0;


SYNTHESIZED_WIRE_20 <= NOT(negDATAandNQ2);



SYNTHESIZED_WIRE_18 <= NOT(NQ1 AND DATA);


NQ1 <= NOT(Q1);



SYNTHESIZED_WIRE_17 <= NOT(Q1 OR NQ2);


SYNTHESIZED_WIRE_16 <= NOT(Q2 OR NQ1 OR Q0);


SYNTHESIZED_WIRE_21 <= Q2 AND Q1;


LOCK <= NOT(NQ0 AND SYNTHESIZED_WIRE_21);


ALARM <= NOT(NQ2 OR NQ1 OR NQ0);


NQ0 <= NOT(Q0);



END bdf_type;